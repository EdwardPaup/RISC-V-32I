import risc_v_32i::*;